
`timescale 1ns/1ns

module test;

reg PCLK,PRESETn,transfer,READ_WRITE;
reg [7:0]apb_write_paddr;
reg [7:0]apb_write_data;
reg [7:0]apb_read_paddr;
wire [7:0]apb_read_data_out;
wire PSLVERR;
reg [7:0]data,expected;

reg [7:0]mem[0:255];

APB_Protocol protocolx(  PCLK,
	                       PRESETn,
		                     transfer,
		                     READ_WRITE,
                         apb_write_paddr,
		                     apb_write_data,
		                     apb_read_paddr,
		                     PSLVERR, 
                         apb_read_data_out);
                         
integer i,j;

initial
begin
  PCLK <= 0;
  forever #5 PCLK = ~PCLK;
end


initial $readmemh("check.mem",mem); 
initial
begin
  PRESETn<=0; transfer<=0; READ_WRITE =0;
  @(posedge PCLK)      PRESETn = 1;                                     //no write address available but request for write operation
  @(posedge PCLK)      transfer = 1;
  repeat(2) @(posedge PCLK);
  @(negedge PCLK)      Write_slave;        // write operation
                               
  repeat(2) @(posedge PCLK);    apb_write_paddr = 8'd22; apb_write_data = 8'd35;
  repeat(2) @(posedge PCLK);
  @(posedge PCLK)     READ_WRITE =1; PRESETn<=0; transfer<=0; 
  @(posedge PCLK)     PRESETn = 1;
  repeat(3) @(posedge PCLK)     transfer = 1;                             // no read address available but request for read operation
  repeat(2) @(posedge PCLK)     Read_slave;                             //read operation

  repeat(3) @(posedge PCLK);   apb_read_paddr = 8'd22;                 //data not inserted in write operation but requested for read operation
  repeat(4) @(posedge PCLK);
  $finish;
end


task Write_slave;
begin
  transfer = 1;
  for (i = 0; i < 8; i = i + 1)
  begin
    repeat(2) @(negedge PCLK)
    begin
      data = i;
      apb_write_data = 2*i;
      apb_write_paddr =  data;
    end
  end
 end 
endtask


 
task Read_slave;
begin
  for (j = 0; j < 8; j = j + 1)
  begin
    repeat(2) @(negedge PCLK)
    begin
      data = j;
      apb_read_paddr =  data;
    end
  end
 end 
endtask


 

  initial
   begin
    $dumpfile("apbWaveform.vcd");
    $dumpvars;
   end

 endmodule
 
 
